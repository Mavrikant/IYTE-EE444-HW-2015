magic
tech scmos
timestamp 1460743457
<< polysilicon >>
rect -20 17 -18 19
rect -12 17 -10 19
rect -4 17 -2 19
rect 4 17 6 19
rect 12 17 14 19
rect 20 17 22 20
rect 28 17 30 20
rect 36 17 38 20
rect -20 10 -18 13
rect -12 10 -10 13
rect -4 10 -2 13
rect 4 10 6 13
rect 12 10 14 13
rect 20 10 22 13
rect 28 10 30 13
rect 36 10 38 13
<< ndiffusion >>
rect -21 13 -20 17
rect -18 13 -17 17
rect -13 13 -12 17
rect -10 13 -9 17
rect -5 13 -4 17
rect -2 13 -1 17
rect 3 13 4 17
rect 6 13 7 17
rect 11 13 12 17
rect 14 13 15 17
rect 19 13 20 17
rect 22 13 23 17
rect 27 13 28 17
rect 30 13 31 17
rect 35 13 36 17
rect 38 13 63 17
<< ntransistor >>
rect -20 13 -18 17
rect -12 13 -10 17
rect -4 13 -2 17
rect 4 13 6 17
rect 12 13 14 17
rect 20 13 22 17
rect 28 13 30 17
rect 36 13 38 17
<< ndcontact >>
rect -25 13 -21 17
rect -17 13 -13 17
rect -9 13 -5 17
rect -1 13 3 17
rect 7 13 11 17
rect 15 13 19 17
rect 23 13 27 17
rect 31 13 35 17
<< end >>
