magic
tech scmos
timestamp 1460379621
<< nwell >>
rect -16 30 0 53
<< polysilicon >>
rect -9 43 -7 45
rect -9 21 -7 31
rect -9 13 -7 15
<< ndiffusion >>
rect -15 20 -9 21
rect -15 16 -14 20
rect -10 16 -9 20
rect -15 15 -9 16
rect -7 20 -1 21
rect -7 16 -6 20
rect -2 16 -1 20
rect -7 15 -1 16
<< pdiffusion >>
rect -15 42 -9 43
rect -15 32 -14 42
rect -10 32 -9 42
rect -15 31 -9 32
rect -7 42 -1 43
rect -7 32 -6 42
rect -2 32 -1 42
rect -7 31 -1 32
<< metal1 >>
rect -16 52 0 53
rect -16 48 -15 52
rect -11 48 -5 52
rect -1 48 0 52
rect -16 47 0 48
rect -14 42 -10 47
rect -6 28 -2 32
rect -16 24 -13 28
rect -6 24 0 28
rect -6 20 -2 24
rect -14 11 -10 16
rect -16 10 0 11
rect -16 6 -15 10
rect -11 6 -5 10
rect -1 6 0 10
rect -16 5 0 6
<< ntransistor >>
rect -9 15 -7 21
<< ptransistor >>
rect -9 31 -7 43
<< polycontact >>
rect -13 24 -9 28
<< ndcontact >>
rect -14 16 -10 20
rect -6 16 -2 20
<< pdcontact >>
rect -14 32 -10 42
rect -6 32 -2 42
<< psubstratepcontact >>
rect -15 6 -11 10
rect -5 6 -1 10
<< nsubstratencontact >>
rect -15 48 -11 52
rect -5 48 -1 52
<< labels >>
rlabel metal1 -8 8 -8 8 1 gnd
rlabel metal1 -8 50 -8 50 5 vcc
rlabel metal1 -15 26 -15 26 3 vin
rlabel metal1 -2 26 -2 26 7 vout
<< end >>
