magic
tech scmos
timestamp 1465466653
<< nwell >>
rect 28 26 464 76
<< polysilicon >>
rect 34 57 36 59
rect 42 57 44 59
rect 83 35 86 39
rect 463 35 465 39
rect 34 25 36 27
rect 42 25 44 27
rect 79 25 83 35
rect 34 23 44 25
rect 50 23 173 25
rect 38 20 40 23
rect 34 11 36 13
rect 42 11 44 13
rect 34 1 36 5
rect 42 1 44 5
rect 50 -11 52 23
rect 171 -11 173 23
rect 182 23 463 25
rect 182 -7 184 23
rect 182 -9 214 -7
rect 50 -13 173 -11
rect 26 -17 35 -15
rect 44 -17 174 -15
rect 202 -17 204 -15
rect 212 -28 214 -9
rect 461 -28 463 23
rect 212 -30 463 -28
<< capacitor >>
rect 52 18 166 23
rect 52 -11 171 18
rect 189 18 461 23
rect 184 -7 461 18
rect 214 -28 461 -7
<< ndiffusion >>
rect 33 5 34 11
rect 36 5 37 11
rect 41 5 42 11
rect 44 5 45 11
rect 35 -15 44 -14
rect 181 -14 202 -10
rect 174 -15 202 -14
rect 35 -18 44 -17
rect 174 -18 202 -17
<< pdiffusion >>
rect 33 27 34 57
rect 36 27 37 57
rect 41 27 42 57
rect 44 27 45 57
rect 93 40 463 47
rect 86 39 463 40
rect 86 34 463 35
rect 86 27 174 34
rect 181 27 463 34
<< metal1 >>
rect 37 74 41 77
rect 37 67 41 70
rect 37 63 93 67
rect 37 57 41 63
rect 86 47 93 63
rect 49 35 79 39
rect 29 20 33 27
rect 29 16 37 20
rect 29 11 33 16
rect 45 11 49 27
rect 174 23 181 27
rect 171 18 184 23
rect 189 18 478 23
rect 37 -10 41 5
rect 174 -10 181 18
rect 44 -22 174 -18
rect 35 -34 44 -22
rect 163 -30 177 -26
rect 189 -30 208 -26
<< ntransistor >>
rect 34 5 36 11
rect 42 5 44 11
rect 35 -17 44 -15
rect 174 -17 202 -15
<< ptransistor >>
rect 34 27 36 57
rect 42 27 44 57
rect 86 35 463 39
<< polycontact >>
rect 79 35 83 39
rect 37 16 41 20
rect 208 -30 212 -26
<< ndcontact >>
rect 29 5 33 11
rect 37 5 41 11
rect 45 5 49 11
rect 35 -14 44 -10
rect 174 -14 181 -10
rect 35 -22 44 -18
rect 174 -22 202 -18
<< pdcontact >>
rect 29 27 33 57
rect 37 27 41 57
rect 45 27 49 57
rect 86 40 93 47
rect 174 27 181 34
<< capcontact >>
rect 166 18 171 23
rect 184 18 189 23
<< psubstratepcontact >>
rect 177 -30 189 -26
<< nsubstratencontact >>
rect 37 70 41 74
<< labels >>
rlabel metal1 472 20 472 20 1 Vout
rlabel metal1 203 -28 203 -28 1 gnd
rlabel polysilicon 35 2 35 2 1 input1
rlabel metal1 38 2 38 2 1 alt
rlabel polysilicon 43 2 43 2 1 input2
rlabel metal1 31 18 31 18 1 orta
rlabel metal1 39 76 39 76 5 vdd
rlabel metal1 52 36 52 36 1 orta2
rlabel metal1 39 -32 39 -32 1 vss
rlabel polysilicon 28 -16 28 -16 3 Vbias
<< end >>
