magic
tech scmos
timestamp 1460911845
<< nwell >>
rect -42 45 84 71
<< polysilicon >>
rect -36 54 -34 56
rect -20 54 -18 56
rect -12 54 -10 56
rect -4 54 -2 56
rect 4 54 6 56
rect 12 54 14 56
rect 20 54 22 56
rect 28 54 30 56
rect 36 54 38 56
rect 44 54 46 56
rect 52 54 54 56
rect 60 54 62 56
rect 68 54 70 56
rect 76 54 78 57
rect -36 33 -34 46
rect -36 27 -34 29
rect -20 17 -18 46
rect -12 17 -10 46
rect -4 17 -2 46
rect 4 17 6 46
rect 12 17 14 46
rect 20 17 22 46
rect 28 17 30 46
rect 36 17 38 46
rect 44 40 46 46
rect 44 17 46 36
rect 52 17 54 46
rect 60 17 62 46
rect 68 17 70 46
rect 76 40 78 46
rect 77 36 78 40
rect 76 17 78 36
rect -20 10 -18 13
rect -12 10 -10 13
rect -4 10 -2 13
rect 4 10 6 13
rect 12 10 14 13
rect 20 10 22 13
rect 28 10 30 13
rect 36 10 38 13
rect 44 11 46 13
rect 52 10 54 13
rect 60 10 62 13
rect 68 10 70 13
rect 76 11 78 13
<< ndiffusion >>
rect -37 29 -36 33
rect -34 29 -33 33
rect -21 13 -20 17
rect -18 13 -17 17
rect -13 13 -12 17
rect -10 13 -9 17
rect -5 13 -4 17
rect -2 13 -1 17
rect 3 13 4 17
rect 6 13 12 17
rect 14 13 15 17
rect 19 13 20 17
rect 22 13 23 17
rect 27 13 28 17
rect 30 13 31 17
rect 35 13 36 17
rect 38 13 39 17
rect 43 13 44 17
rect 46 13 47 17
rect 51 13 52 17
rect 54 13 60 17
rect 62 13 68 17
rect 70 13 71 17
rect 75 13 76 17
rect 78 13 79 17
<< pdiffusion >>
rect -37 46 -36 54
rect -34 46 -33 54
rect -21 46 -20 54
rect -18 46 -17 54
rect -13 46 -12 54
rect -10 46 -9 54
rect -5 46 -4 54
rect -2 46 -1 54
rect 3 46 4 54
rect 6 46 12 54
rect 14 46 15 54
rect 19 46 20 54
rect 22 46 23 54
rect 27 46 28 54
rect 30 46 31 54
rect 35 46 36 54
rect 38 46 39 54
rect 43 46 44 54
rect 46 46 47 54
rect 51 46 52 54
rect 54 46 60 54
rect 62 46 68 54
rect 70 46 71 54
rect 75 46 76 54
rect 78 46 79 54
<< metal1 >>
rect 15 70 19 80
rect -29 66 15 70
rect 19 66 71 70
rect -33 54 -29 66
rect -25 54 -21 58
rect -17 54 -13 66
rect -9 54 -5 58
rect 15 54 19 66
rect 23 54 27 58
rect 31 54 35 66
rect 39 54 43 58
rect 71 54 75 66
rect 51 46 59 54
rect 79 54 83 80
rect -41 41 -38 46
rect -46 37 -38 41
rect -1 40 3 46
rect 55 40 59 46
rect -41 33 -38 37
rect -30 36 -1 40
rect 3 36 43 40
rect 59 36 73 40
rect -29 29 75 33
rect -33 -31 -29 29
rect -25 17 -21 21
rect -17 17 -13 29
rect -9 17 -5 21
rect -1 17 3 21
rect 15 17 19 29
rect 23 17 27 21
rect 31 17 35 29
rect 39 17 43 21
rect 55 17 59 21
rect 51 13 59 17
rect 71 17 75 29
rect 80 17 83 46
rect 86 37 94 41
rect 86 10 90 37
rect -21 -6 -17 6
rect -13 2 -9 6
rect -5 2 -1 6
rect 3 -6 7 6
rect 11 2 15 6
rect 19 2 23 6
rect 27 -6 31 6
rect 35 2 39 6
rect 51 -6 55 6
rect -21 -10 55 -6
rect -21 -31 -17 -10
rect 59 -14 63 6
rect -9 -18 11 -14
rect 15 -18 35 -14
rect 39 -18 63 -14
rect 71 6 90 10
rect -13 -31 -9 -18
rect 67 -22 71 6
rect -1 -26 19 -22
rect 23 -26 71 -22
<< metal2 >>
rect -21 58 -9 62
rect 27 58 39 62
rect -1 25 3 36
rect 55 25 59 36
rect -21 21 -9 25
rect 27 21 39 25
rect -13 -14 -9 -2
rect -5 -22 -1 -2
rect 11 -14 15 -2
rect 19 -22 23 -2
rect 35 -14 39 -2
<< ntransistor >>
rect -36 29 -34 33
rect -20 13 -18 17
rect -12 13 -10 17
rect -4 13 -2 17
rect 4 13 6 17
rect 12 13 14 17
rect 20 13 22 17
rect 28 13 30 17
rect 36 13 38 17
rect 44 13 46 17
rect 52 13 54 17
rect 60 13 62 17
rect 68 13 70 17
rect 76 13 78 17
<< ptransistor >>
rect -36 46 -34 54
rect -20 46 -18 54
rect -12 46 -10 54
rect -4 46 -2 54
rect 4 46 6 54
rect 12 46 14 54
rect 20 46 22 54
rect 28 46 30 54
rect 36 46 38 54
rect 44 46 46 54
rect 52 46 54 54
rect 60 46 62 54
rect 68 46 70 54
rect 76 46 78 54
<< polycontact >>
rect -34 36 -30 40
rect 43 36 47 40
rect 73 36 77 40
rect -21 6 -17 10
rect -13 6 -9 10
rect -5 6 -1 10
rect 3 6 7 10
rect 11 6 15 10
rect 19 6 23 10
rect 27 6 31 10
rect 35 6 39 10
rect 51 6 55 10
rect 59 6 63 10
rect 67 6 71 10
<< ndcontact >>
rect -41 29 -37 33
rect -33 29 -29 33
rect -25 13 -21 17
rect -17 13 -13 17
rect -9 13 -5 17
rect -1 13 3 17
rect 15 13 19 17
rect 23 13 27 17
rect 31 13 35 17
rect 39 13 43 17
rect 47 13 51 17
rect 71 13 75 17
rect 79 13 83 17
<< pdcontact >>
rect -41 46 -37 54
rect -33 46 -29 54
rect -25 46 -21 54
rect -17 46 -13 54
rect -9 46 -5 54
rect -1 46 3 54
rect 15 46 19 54
rect 23 46 27 54
rect 31 46 35 54
rect 39 46 43 54
rect 47 46 51 54
rect 71 46 75 54
rect 79 46 83 54
<< m2contact >>
rect -25 58 -21 62
rect -9 58 -5 62
rect 23 58 27 62
rect 39 58 43 62
rect -1 36 3 40
rect 55 36 59 40
rect -25 21 -21 25
rect -9 21 -5 25
rect -1 21 3 25
rect 23 21 27 25
rect 39 21 43 25
rect 55 21 59 25
rect -13 -2 -9 2
rect -5 -2 -1 2
rect 11 -2 15 2
rect 19 -2 23 2
rect 35 -2 39 2
rect -13 -18 -9 -14
rect 11 -18 15 -14
rect 35 -18 39 -14
rect -5 -26 -1 -22
rect 19 -26 23 -22
<< nsubstratencontact >>
rect -33 66 -29 70
rect 15 66 19 70
rect 71 66 75 70
<< labels >>
rlabel metal1 -45 39 -45 39 3 Cout
rlabel metal1 81 79 81 79 6 Sum
rlabel metal1 -31 -29 -31 -29 1 Gnd
rlabel metal1 -19 -29 -19 -29 1 A
rlabel metal1 -11 -29 -11 -29 1 B
rlabel metal1 93 39 93 39 7 Cin
rlabel metal1 17 79 17 79 5 Vdd
<< end >>
