magic
tech scmos
timestamp 1460748030
<< polysilicon >>
rect -20 17 -18 46
rect -12 17 -10 44
rect -4 17 -2 45
rect 4 17 6 38
rect 12 17 14 41
rect 20 17 22 45
rect 28 17 30 46
rect 36 17 38 44
rect 44 17 46 45
rect 52 17 54 45
rect 60 17 62 47
rect 68 17 70 47
rect 76 17 78 48
rect -20 10 -18 13
rect -12 10 -10 13
rect -4 10 -2 13
rect 4 10 6 13
rect 12 10 14 13
rect 20 10 22 13
rect 28 10 30 13
rect 36 10 38 13
rect 44 10 46 13
rect 52 10 54 13
rect 60 10 62 13
rect 68 10 70 13
rect 76 10 78 13
<< ndiffusion >>
rect -21 13 -20 17
rect -18 13 -17 17
rect -13 13 -12 17
rect -10 13 -9 17
rect -5 13 -4 17
rect -2 13 -1 17
rect 3 13 4 17
rect 6 13 7 17
rect 11 13 12 17
rect 14 13 15 17
rect 19 13 20 17
rect 22 13 23 17
rect 27 13 28 17
rect 30 13 31 17
rect 35 13 36 17
rect 38 13 39 17
rect 43 13 44 17
rect 46 13 47 17
rect 51 13 52 17
rect 54 13 55 17
rect 59 13 60 17
rect 62 13 63 17
rect 67 13 68 17
rect 70 13 71 17
rect 75 13 76 17
rect 78 13 79 17
<< metal1 >>
rect -17 29 55 33
rect 79 29 83 32
rect -25 17 -21 21
rect -17 17 -13 29
rect 79 25 104 29
rect 63 21 112 25
rect -9 17 -5 21
rect 79 17 83 21
rect -21 -6 -17 6
rect -13 2 -9 6
rect -5 2 -1 6
rect 3 -6 7 6
rect 11 2 15 6
rect 19 2 23 6
rect 27 -6 31 6
rect 35 2 39 6
rect 43 2 47 6
rect 51 2 55 6
rect 59 2 63 6
rect 67 2 71 6
rect 75 -6 79 6
rect -28 -10 80 -6
rect -28 -18 -13 -14
rect -9 -18 11 -14
rect 15 -18 35 -14
rect 39 -18 67 -14
rect 71 -18 80 -14
rect -28 -26 -5 -22
rect -1 -26 19 -22
rect 23 -26 59 -22
rect 63 -26 80 -22
<< metal2 >>
rect -21 21 -9 25
rect -13 -14 -9 -2
rect -5 -22 -1 -2
rect 11 -14 15 -2
rect 19 -22 23 -2
rect 35 -14 39 -2
rect 59 -22 63 -2
rect 67 -14 71 -2
<< ntransistor >>
rect -20 13 -18 17
rect -12 13 -10 17
rect -4 13 -2 17
rect 4 13 6 17
rect 12 13 14 17
rect 20 13 22 17
rect 28 13 30 17
rect 36 13 38 17
rect 44 13 46 17
rect 52 13 54 17
rect 60 13 62 17
rect 68 13 70 17
rect 76 13 78 17
<< polycontact >>
rect -21 6 -17 10
rect -13 6 -9 10
rect -5 6 -1 10
rect 3 6 7 10
rect 11 6 15 10
rect 19 6 23 10
rect 27 6 31 10
rect 35 6 39 10
rect 43 6 47 10
rect 51 6 55 10
rect 59 6 63 10
rect 67 6 71 10
rect 75 6 79 10
<< ndcontact >>
rect -25 13 -21 17
rect -17 13 -13 17
rect -9 13 -5 17
rect -1 13 3 17
rect 7 13 11 17
rect 15 13 19 17
rect 23 13 27 17
rect 31 13 35 17
rect 39 13 43 17
rect 47 13 51 17
rect 55 13 59 17
rect 63 13 67 17
rect 71 13 75 17
rect 79 13 83 17
<< m2contact >>
rect -25 21 -21 25
rect -9 21 -5 25
rect -13 -2 -9 2
rect -5 -2 -1 2
rect 11 -2 15 2
rect 19 -2 23 2
rect 35 -2 39 2
rect 59 -2 63 2
rect 67 -2 71 2
rect -13 -18 -9 -14
rect 11 -18 15 -14
rect 35 -18 39 -14
rect 67 -18 71 -14
rect -5 -26 -1 -22
rect 19 -26 23 -22
rect 59 -26 63 -22
<< end >>
