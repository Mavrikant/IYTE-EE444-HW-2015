magic
tech scmos
timestamp 1461970242
<< nwell >>
rect 147 56 261 79
<< polysilicon >>
rect 170 69 225 71
rect 157 65 159 67
rect 167 65 169 68
rect 177 65 179 67
rect 187 65 189 67
rect 205 65 207 69
rect 223 65 225 69
rect 233 65 235 68
rect 243 65 245 67
rect 253 65 255 67
rect 157 52 159 57
rect 167 55 169 57
rect 177 53 179 57
rect 157 50 169 52
rect 157 45 159 47
rect 167 45 169 50
rect 177 49 178 53
rect 177 45 179 49
rect 187 45 189 57
rect 205 45 207 57
rect 223 52 225 57
rect 233 55 235 57
rect 243 53 245 57
rect 223 50 235 52
rect 223 45 225 47
rect 233 45 235 50
rect 243 49 244 53
rect 243 45 245 49
rect 253 45 255 57
rect 157 38 159 41
rect 158 34 159 38
rect 167 31 169 41
rect 177 39 179 41
rect 187 38 189 41
rect 205 39 207 41
rect 187 34 188 38
rect 223 32 225 41
rect 233 39 235 41
rect 243 39 245 41
rect 253 38 255 41
rect 253 34 257 38
rect 199 31 203 32
rect 167 29 217 31
rect 221 28 225 32
<< ndiffusion >>
rect 155 41 157 45
rect 159 41 161 45
rect 165 41 167 45
rect 169 41 171 45
rect 175 41 177 45
rect 179 41 181 45
rect 185 41 187 45
rect 189 41 191 45
rect 203 41 205 45
rect 207 41 209 45
rect 221 41 223 45
rect 225 41 227 45
rect 231 41 233 45
rect 235 41 237 45
rect 241 41 243 45
rect 245 41 247 45
rect 251 41 253 45
rect 255 41 257 45
<< pdiffusion >>
rect 155 57 157 65
rect 159 57 161 65
rect 165 57 167 65
rect 169 57 171 65
rect 175 57 177 65
rect 179 57 181 65
rect 185 57 187 65
rect 189 57 191 65
rect 203 57 205 65
rect 207 57 209 65
rect 221 57 223 65
rect 225 57 227 65
rect 231 57 233 65
rect 235 57 237 65
rect 241 57 243 65
rect 245 57 247 65
rect 251 57 253 65
rect 255 57 257 65
<< metal1 >>
rect 137 75 151 79
rect 155 75 169 79
rect 173 75 195 79
rect 199 75 217 79
rect 221 75 235 79
rect 239 75 257 79
rect 137 68 149 72
rect 153 68 166 72
rect 181 65 185 75
rect 209 65 213 75
rect 236 68 237 72
rect 247 65 251 75
rect 151 53 155 57
rect 137 49 155 53
rect 151 45 155 49
rect 161 45 165 57
rect 171 53 175 57
rect 191 53 195 57
rect 182 49 195 53
rect 171 45 175 49
rect 191 45 195 49
rect 199 45 203 57
rect 217 53 221 57
rect 213 49 221 53
rect 217 45 221 49
rect 153 34 154 38
rect 161 33 165 41
rect 181 40 185 41
rect 188 33 192 34
rect 161 30 192 33
rect 199 36 203 41
rect 227 45 231 57
rect 237 53 241 57
rect 257 53 261 57
rect 248 49 261 53
rect 237 45 241 49
rect 257 45 261 49
rect 209 40 213 41
rect 217 32 221 34
rect 137 26 147 30
rect 151 26 154 30
rect 227 33 231 41
rect 247 40 251 41
rect 257 33 261 34
rect 227 29 261 33
<< metal2 >>
rect 149 38 153 68
rect 217 68 237 72
rect 175 49 209 53
rect 181 30 185 36
rect 209 30 213 36
rect 217 38 221 68
rect 241 49 265 53
rect 247 30 251 36
rect 158 26 261 30
<< ntransistor >>
rect 157 41 159 45
rect 167 41 169 45
rect 177 41 179 45
rect 187 41 189 45
rect 205 41 207 45
rect 223 41 225 45
rect 233 41 235 45
rect 243 41 245 45
rect 253 41 255 45
<< ptransistor >>
rect 157 57 159 65
rect 167 57 169 65
rect 177 57 179 65
rect 187 57 189 65
rect 205 57 207 65
rect 223 57 225 65
rect 233 57 235 65
rect 243 57 245 65
rect 253 57 255 65
<< polycontact >>
rect 166 68 170 72
rect 232 68 236 72
rect 178 49 182 53
rect 244 49 248 53
rect 154 34 158 38
rect 188 34 192 38
rect 199 32 203 36
rect 257 34 261 38
rect 217 28 221 32
<< ndcontact >>
rect 151 41 155 45
rect 161 41 165 45
rect 171 41 175 45
rect 181 41 185 45
rect 191 41 195 45
rect 199 41 203 45
rect 209 41 213 45
rect 217 41 221 45
rect 227 41 231 45
rect 237 41 241 45
rect 247 41 251 45
rect 257 41 261 45
<< pdcontact >>
rect 151 57 155 65
rect 161 57 165 65
rect 171 57 175 65
rect 181 57 185 65
rect 191 57 195 65
rect 199 57 203 65
rect 209 57 213 65
rect 217 57 221 65
rect 227 57 231 65
rect 237 57 241 65
rect 247 57 251 65
rect 257 57 261 65
<< m2contact >>
rect 149 68 153 72
rect 237 68 241 72
rect 171 49 175 53
rect 209 49 213 53
rect 149 34 153 38
rect 181 36 185 40
rect 237 49 241 53
rect 209 36 213 40
rect 217 34 221 38
rect 154 26 158 30
rect 247 36 251 40
<< psubstratepcontact >>
rect 147 26 151 30
<< nsubstratencontact >>
rect 151 75 155 79
rect 169 75 173 79
rect 195 75 199 79
rect 217 75 221 79
rect 235 75 239 79
rect 257 75 261 79
<< labels >>
rlabel metal1 138 77 138 77 4 Vdd
rlabel metal1 138 70 138 70 3 Clk
rlabel metal1 138 28 138 28 2 Gnd
rlabel metal1 148 51 148 51 3 D
rlabel metal1 214 51 214 51 7 Q1
rlabel metal2 263 51 263 51 7 Q2
<< end >>
