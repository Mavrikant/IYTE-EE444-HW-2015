magic
tech scmos
timestamp 1460746148
<< polysilicon >>
rect -20 43 -18 47
rect -12 43 -10 47
rect -4 43 -2 47
rect 4 43 6 47
rect 12 43 14 47
rect 20 43 22 47
rect 28 43 30 47
rect 36 43 38 47
rect 44 43 46 47
rect 52 43 54 47
rect 60 43 62 47
rect 68 43 70 47
rect 76 43 78 47
rect -20 17 -18 35
rect -12 17 -10 35
rect -4 17 -2 35
rect 4 17 6 35
rect 12 17 14 35
rect 20 17 22 35
rect 28 17 30 35
rect 36 17 38 35
rect 44 17 46 35
rect 52 17 54 35
rect 60 17 62 35
rect 68 17 70 35
rect 76 17 78 35
rect -20 10 -18 13
rect -12 10 -10 13
rect -4 10 -2 13
rect 4 10 6 13
rect 12 10 14 13
rect 20 10 22 13
rect 28 10 30 13
rect 36 10 38 13
rect 44 10 46 13
rect 52 10 54 13
rect 60 10 62 13
rect 68 10 70 13
rect 76 10 78 13
<< ndiffusion >>
rect -21 13 -20 17
rect -18 13 -17 17
rect -13 13 -12 17
rect -10 13 -9 17
rect -5 13 -4 17
rect -2 13 -1 17
rect 3 13 4 17
rect 6 13 7 17
rect 11 13 12 17
rect 14 13 15 17
rect 19 13 20 17
rect 22 13 23 17
rect 27 13 28 17
rect 30 13 31 17
rect 35 13 36 17
rect 38 13 39 17
rect 43 13 44 17
rect 46 13 47 17
rect 51 13 52 17
rect 54 13 55 17
rect 59 13 60 17
rect 62 13 63 17
rect 67 13 68 17
rect 70 13 71 17
rect 75 13 76 17
rect 78 13 79 17
<< pdiffusion >>
rect -21 35 -20 43
rect -18 35 -17 43
rect -13 35 -12 43
rect -10 35 -9 43
rect -5 35 -4 43
rect -2 35 -1 43
rect 3 35 4 43
rect 6 35 7 43
rect 11 35 12 43
rect 14 35 15 43
rect 19 35 20 43
rect 22 35 23 43
rect 27 35 28 43
rect 30 35 31 43
rect 35 35 36 43
rect 38 35 39 43
rect 43 35 44 43
rect 46 35 47 43
rect 51 35 52 43
rect 54 35 55 43
rect 59 35 60 43
rect 62 35 63 43
rect 67 35 68 43
rect 70 35 71 43
rect 75 35 76 43
rect 78 35 79 43
<< metal1 >>
rect -41 35 -25 43
rect 79 29 83 35
rect 79 25 104 29
rect 79 17 83 25
rect -38 13 -25 17
rect -21 -6 -17 6
rect -13 2 -9 6
rect -5 2 -1 6
rect 3 -6 7 6
rect 11 2 15 6
rect 19 2 23 6
rect 27 -6 31 6
rect 35 2 39 6
rect 43 2 47 6
rect 51 2 55 6
rect 59 2 63 6
rect 67 2 71 6
rect 75 -6 79 6
rect -28 -10 80 -6
rect -28 -18 -13 -14
rect -9 -18 11 -14
rect 15 -18 35 -14
rect 39 -18 67 -14
rect 71 -18 80 -14
rect -28 -26 -5 -22
rect -1 -26 19 -22
rect 23 -26 59 -22
rect 63 -26 80 -22
<< metal2 >>
rect -13 -14 -9 -2
rect -5 -22 -1 -2
rect 11 -14 15 -2
rect 19 -22 23 -2
rect 35 -14 39 -2
rect 59 -22 63 -2
rect 67 -14 71 -2
<< ntransistor >>
rect -20 13 -18 17
rect -12 13 -10 17
rect -4 13 -2 17
rect 4 13 6 17
rect 12 13 14 17
rect 20 13 22 17
rect 28 13 30 17
rect 36 13 38 17
rect 44 13 46 17
rect 52 13 54 17
rect 60 13 62 17
rect 68 13 70 17
rect 76 13 78 17
<< ptransistor >>
rect -20 35 -18 43
rect -12 35 -10 43
rect -4 35 -2 43
rect 4 35 6 43
rect 12 35 14 43
rect 20 35 22 43
rect 28 35 30 43
rect 36 35 38 43
rect 44 35 46 43
rect 52 35 54 43
rect 60 35 62 43
rect 68 35 70 43
rect 76 35 78 43
<< polycontact >>
rect -21 6 -17 10
rect -13 6 -9 10
rect -5 6 -1 10
rect 3 6 7 10
rect 11 6 15 10
rect 19 6 23 10
rect 27 6 31 10
rect 35 6 39 10
rect 43 6 47 10
rect 51 6 55 10
rect 59 6 63 10
rect 67 6 71 10
rect 75 6 79 10
<< ndcontact >>
rect -25 13 -21 17
rect -17 13 -13 17
rect -9 13 -5 17
rect -1 13 3 17
rect 7 13 11 17
rect 15 13 19 17
rect 23 13 27 17
rect 31 13 35 17
rect 39 13 43 17
rect 47 13 51 17
rect 55 13 59 17
rect 63 13 67 17
rect 71 13 75 17
rect 79 13 83 17
<< pdcontact >>
rect -25 35 -21 43
rect -17 35 -13 43
rect -9 35 -5 43
rect -1 35 3 43
rect 7 35 11 43
rect 15 35 19 43
rect 23 35 27 43
rect 31 35 35 43
rect 39 35 43 43
rect 47 35 51 43
rect 55 35 59 43
rect 63 35 67 43
rect 71 35 75 43
rect 79 35 83 43
<< m2contact >>
rect -13 -2 -9 2
rect -5 -2 -1 2
rect 11 -2 15 2
rect 19 -2 23 2
rect 35 -2 39 2
rect 59 -2 63 2
rect 67 -2 71 2
rect -13 -18 -9 -14
rect 11 -18 15 -14
rect 35 -18 39 -14
rect 67 -18 71 -14
rect -5 -26 -1 -22
rect 19 -26 23 -22
rect 59 -26 63 -22
<< end >>
