* M. Serdar Karaman
* 190206038

.model nfet NMOS
.model pfet PMOS

M1000 vout vin vcc vcc pfet w=12 l=2
+  ad=72 pd=36 as=72 ps=36

M1001 vout vin gnd Gnd nfet w=6 l=2
+  ad=36 pd=24 as=36 ps=24

* SPICE language is case insensitive, ignore this Gnd-gnd cap.
C0 gnd Gnd 3.8fF 
C1 vout Gnd 2.1fF
C2 vin Gnd 4.9fF

V1 vin Gnd PULSE(0 5 0 1f 1f .125n .25n )
V2 vcc Gnd 5

.tran 10000n 1ns
.end
